interface er_simple_clk_reset_if();
   bit clk,nreset;
endinterface // er_simple_clk_reset_if
