// *************************************************************************************
// Copyright 2014 Mentor Graphics Corporation
// All Rights Reserved
//
// THIS WORK CONTAINS TRADE SECRET AND PROPRIETARY INFORMATION WHICH IS THE PROPERTY OF
// MENTOR GRAPHICS CORPORATION OR ITS LICENSORS AND IS SUBJECT TO LICENSE TERMS
//
// bugs, enhancement requests to: avidan_efody@mentor.com
// *************************************************************************************

interface sli_clk_reset_if();
   bit clk,nreset;
endinterface // sli_clk_reset_if
