interface er_tap_1500_if(input WRCK,WRSTN);

// Naming as of standard
bit WSI, WSO, SelectWIR, CaptureWR, ShiftWR,UpdateWR;
// Optional
bit TransferDR;



endinterface
