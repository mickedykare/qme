//----------------------------------------------------------------------
//                   Mentor Graphics Corporation
//----------------------------------------------------------------------
// Project         : generic_reg_bus_agent
// Unit            : ra_example_tb_pkg
// File            : ra_example_tb_pkg.svh
//----------------------------------------------------------------------
// Created by      : mikaela
// Creation Date   : 2014/06/05
//----------------------------------------------------------------------
// Title: 
//
// Summary:
//
// Description:
//
//----------------------------------------------------------------------

//----------------------------------------------------------------------
// ra_example_tb_pkg
//----------------------------------------------------------------------
package ra_example_tb_pkg;

  `include "uvm_macros.svh"  
   import uvm_pkg::*;
   import example_block_regs_pkg::*;
   import apb3_uvm_reg_pkg::*;
   import mvc_pkg::*;
   import mgc_apb3_v1_0_pkg::*; 
   import sli_clk_reset_pkg::*;
   

  `include "ra_example_tb_env.svh"
  `include "ra_example_base_test.svh"
   
   
   
   
endpackage: ra_example_tb_pkg

