../src/vhdl/components.vhd
../src/vhdl/qft_lib.vhd
../src/vhdl/pinmux.vhd
../src/vhdl/apb_master_sc.vhd
../src/vhdl/apb_access_arb.vhd
../src/vhdl/apb_master_mc.vhd
../src/vhdl/master_interface.vhd
../src/vhdl/axi4lite_slave.vhd
../src/vhdl/dp_sram.vhd
../src/vhdl/dp_fifo.vhd
../src/vhdl/fifos.vhd
../src/vhdl/apb_slave_int.vhd
../src/vhdl/config_status_reg.vhd
../src/vhdl/csr_interface_apb.vhd
../src/vhdl/axi4lite_to_apb4.vhd
